VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_8_8192_scn4m_subm
   CLASS BLOCK ;
   SIZE 1260.5 BY 5799.6 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  282.2 0.0 283.4 1.2 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  304.0 0.0 305.2 1.2 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  325.8 0.0 327.0 1.2 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  347.6 0.0 348.8 1.2 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  369.4 0.0 370.6 1.2 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  391.2 0.0 392.4 1.2 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  413.0 0.0 414.2 1.2 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  434.8 0.0 436.0 1.2 ;
      END
   END din0[7]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  195.0 0.0 196.2 1.2 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  216.8 0.0 218.0 1.2 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  238.6 0.0 239.8 1.2 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  260.4 0.0 261.6 1.2 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 734.2 1.2 735.4 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 756.2 1.2 757.4 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 774.2 1.2 775.4 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 796.2 1.2 797.4 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 814.2 1.2 815.4 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 836.2 1.2 837.4 ;
      END
   END addr0[9]
   PIN addr0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 854.2 1.2 855.4 ;
      END
   END addr0[10]
   PIN addr0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 876.2 1.2 877.4 ;
      END
   END addr0[11]
   PIN addr0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 894.2 1.2 895.4 ;
      END
   END addr0[12]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 258.0 1.2 259.2 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 280.0 1.2 281.2 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 260.0 1.2 261.2 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  345.0 0.0 346.2 1.2 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  457.1 0.0 458.3 1.2 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  565.9 0.0 567.1 1.2 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  674.7 0.0 675.9 1.2 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  783.5 0.0 784.7 1.2 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  892.3 0.0 893.5 1.2 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  1259.3 299.2 1260.5 300.4 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  1259.3 301.2 1260.5 302.4 ;
      END
   END dout0[7]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  0.0 5793.6 1260.5 5799.6 ;
         LAYER metal4 ;
         RECT  1254.5 0.0 1260.5 5799.6 ;
         LAYER metal4 ;
         RECT  0.0 0.0 6.0 5799.6 ;
         LAYER metal3 ;
         RECT  0.0 0.0 1260.5 6.0 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  12.0 12.0 18.0 5787.6 ;
         LAYER metal4 ;
         RECT  1242.5 12.0 1248.5 5787.6 ;
         LAYER metal3 ;
         RECT  12.0 5781.6 1248.5 5787.6 ;
         LAYER metal3 ;
         RECT  12.0 12.0 1248.5 18.0 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  1.4 1.4 1259.1 5798.2 ;
   LAYER  metal2 ;
      RECT  1.4 1.4 1259.1 5798.2 ;
   LAYER  metal3 ;
      RECT  2.4 733.0 1259.1 736.6 ;
      RECT  1.4 736.6 2.4 755.0 ;
      RECT  1.4 758.6 2.4 773.0 ;
      RECT  1.4 776.6 2.4 795.0 ;
      RECT  1.4 798.6 2.4 813.0 ;
      RECT  1.4 816.6 2.4 835.0 ;
      RECT  1.4 838.6 2.4 853.0 ;
      RECT  1.4 856.6 2.4 875.0 ;
      RECT  1.4 878.6 2.4 893.0 ;
      RECT  1.4 282.4 2.4 733.0 ;
      RECT  1.4 262.4 2.4 278.8 ;
      RECT  2.4 298.0 1258.1 301.6 ;
      RECT  2.4 301.6 1258.1 733.0 ;
      RECT  1258.1 303.6 1259.1 733.0 ;
      RECT  1.4 896.6 2.4 5792.4 ;
      RECT  1.4 7.2 2.4 256.8 ;
      RECT  1258.1 7.2 1259.1 298.0 ;
      RECT  2.4 736.6 10.8 5780.4 ;
      RECT  2.4 5780.4 10.8 5788.8 ;
      RECT  2.4 5788.8 10.8 5792.4 ;
      RECT  10.8 736.6 1249.7 5780.4 ;
      RECT  10.8 5788.8 1249.7 5792.4 ;
      RECT  1249.7 736.6 1259.1 5780.4 ;
      RECT  1249.7 5780.4 1259.1 5788.8 ;
      RECT  1249.7 5788.8 1259.1 5792.4 ;
      RECT  2.4 7.2 10.8 10.8 ;
      RECT  2.4 10.8 10.8 19.2 ;
      RECT  2.4 19.2 10.8 298.0 ;
      RECT  10.8 7.2 1249.7 10.8 ;
      RECT  10.8 19.2 1249.7 298.0 ;
      RECT  1249.7 7.2 1258.1 10.8 ;
      RECT  1249.7 10.8 1258.1 19.2 ;
      RECT  1249.7 19.2 1258.1 298.0 ;
   LAYER  metal4 ;
      RECT  279.8 3.6 285.8 5798.2 ;
      RECT  285.8 1.4 301.6 3.6 ;
      RECT  307.6 1.4 323.4 3.6 ;
      RECT  351.2 1.4 367.0 3.6 ;
      RECT  373.0 1.4 388.8 3.6 ;
      RECT  394.8 1.4 410.6 3.6 ;
      RECT  416.6 1.4 432.4 3.6 ;
      RECT  198.6 1.4 214.4 3.6 ;
      RECT  220.4 1.4 236.2 3.6 ;
      RECT  242.2 1.4 258.0 3.6 ;
      RECT  264.0 1.4 279.8 3.6 ;
      RECT  329.4 1.4 342.6 3.6 ;
      RECT  438.4 1.4 454.7 3.6 ;
      RECT  460.7 1.4 563.5 3.6 ;
      RECT  569.5 1.4 672.3 3.6 ;
      RECT  678.3 1.4 781.1 3.6 ;
      RECT  787.1 1.4 889.9 3.6 ;
      RECT  895.9 1.4 1252.1 3.6 ;
      RECT  8.4 1.4 192.6 3.6 ;
      RECT  8.4 3.6 9.6 9.6 ;
      RECT  8.4 9.6 9.6 5790.0 ;
      RECT  8.4 5790.0 9.6 5798.2 ;
      RECT  9.6 3.6 20.4 9.6 ;
      RECT  9.6 5790.0 20.4 5798.2 ;
      RECT  20.4 3.6 279.8 9.6 ;
      RECT  20.4 9.6 279.8 5790.0 ;
      RECT  20.4 5790.0 279.8 5798.2 ;
      RECT  285.8 3.6 1240.1 9.6 ;
      RECT  285.8 9.6 1240.1 5790.0 ;
      RECT  285.8 5790.0 1240.1 5798.2 ;
      RECT  1240.1 3.6 1250.9 9.6 ;
      RECT  1240.1 5790.0 1250.9 5798.2 ;
      RECT  1250.9 3.6 1252.1 9.6 ;
      RECT  1250.9 9.6 1252.1 5790.0 ;
      RECT  1250.9 5790.0 1252.1 5798.2 ;
   END
END    sram_8_8192_scn4m_subm
END    LIBRARY
